simple test for names = ft_getpnames() versus free_pnode(names)

.control
let buf = [ 1 2 3 ]
let buf2=db(mag(buf))
quit
.endc

.end
