simple test for names = ft_getpnames() versus free_pnode(names)

.control
let buf = 0
let buf = buf + 1
quit
.endc

.end
